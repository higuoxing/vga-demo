`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/31/2017 03:10:15 AM
// Design Name: 
// Module Name: cross_hair_handler
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module cross_hair_handler(clk, hsync, vsync, hcnt, vcnt, hcnt_out, vcnt_out);

//    input clk, hsync, vsync, hcnt, vcnt;
//    output hcnt_out, vcnt_out;
    
//    wire clk, hsync, vsync;
//    wire [9:0] hcnt, vcnt;
//    reg [9:0] hcnt_out, vcnt_out;
    
//    always @ (posedge(clk)) begin
        
//        if (vsync) begin
        
//            hcnt_out <= 0;
//            vcnt_out <= 0;
            
//    end
    
//endmodule
